`timescale 1ns / 1ps


module KSadd8(
    input [7:0] a,
    input [7:0] b,
    input cin,
    output [7:0] sum,
    output cout;
    );
endmodule
